module gw_gao(
    \digital_out[7] ,
    \digital_out[6] ,
    \digital_out[5] ,
    \digital_out[4] ,
    \digital_out[3] ,
    \digital_out[2] ,
    \digital_out[1] ,
    \digital_out[0] ,
    \SSD_ADC/accum[7] ,
    \SSD_ADC/accum[6] ,
    \SSD_ADC/accum[5] ,
    \SSD_ADC/accum[4] ,
    \SSD_ADC/accum[3] ,
    \SSD_ADC/accum[2] ,
    \SSD_ADC/accum[1] ,
    \SSD_ADC/accum[0] ,
    \SSD_ADC/accum_rdy ,
    analog_out,
    analog_cmp,
    clk,
    sample_rdy,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \digital_out[7] ;
input \digital_out[6] ;
input \digital_out[5] ;
input \digital_out[4] ;
input \digital_out[3] ;
input \digital_out[2] ;
input \digital_out[1] ;
input \digital_out[0] ;
input \SSD_ADC/accum[7] ;
input \SSD_ADC/accum[6] ;
input \SSD_ADC/accum[5] ;
input \SSD_ADC/accum[4] ;
input \SSD_ADC/accum[3] ;
input \SSD_ADC/accum[2] ;
input \SSD_ADC/accum[1] ;
input \SSD_ADC/accum[0] ;
input \SSD_ADC/accum_rdy ;
input analog_out;
input analog_cmp;
input clk;
input sample_rdy;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \digital_out[7] ;
wire \digital_out[6] ;
wire \digital_out[5] ;
wire \digital_out[4] ;
wire \digital_out[3] ;
wire \digital_out[2] ;
wire \digital_out[1] ;
wire \digital_out[0] ;
wire \SSD_ADC/accum[7] ;
wire \SSD_ADC/accum[6] ;
wire \SSD_ADC/accum[5] ;
wire \SSD_ADC/accum[4] ;
wire \SSD_ADC/accum[3] ;
wire \SSD_ADC/accum[2] ;
wire \SSD_ADC/accum[1] ;
wire \SSD_ADC/accum[0] ;
wire \SSD_ADC/accum_rdy ;
wire analog_out;
wire analog_cmp;
wire clk;
wire sample_rdy;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i({\digital_out[7] ,\digital_out[6] ,\digital_out[5] ,\digital_out[4] ,\digital_out[3] ,\digital_out[2] ,\digital_out[1] ,\digital_out[0] ,\SSD_ADC/accum[7] ,\SSD_ADC/accum[6] ,\SSD_ADC/accum[5] ,\SSD_ADC/accum[4] ,\SSD_ADC/accum[3] ,\SSD_ADC/accum[2] ,\SSD_ADC/accum[1] ,\SSD_ADC/accum[0] ,\SSD_ADC/accum_rdy ,analog_out,analog_cmp,clk,sample_rdy}),
    .trig1_i(sample_rdy),
    .data_i({\digital_out[7] ,\digital_out[6] ,\digital_out[5] ,\digital_out[4] ,\digital_out[3] ,\digital_out[2] ,\digital_out[1] ,\digital_out[0] ,\SSD_ADC/accum[7] ,\SSD_ADC/accum[6] ,\SSD_ADC/accum[5] ,\SSD_ADC/accum[4] ,\SSD_ADC/accum[3] ,\SSD_ADC/accum[2] ,\SSD_ADC/accum[1] ,\SSD_ADC/accum[0] ,\SSD_ADC/accum_rdy ,analog_out,analog_cmp,clk,sample_rdy}),
    .clk_i(clk)
);

endmodule
